
-- Module : divisor
-- Author : folletto
-- Date   : gio, 1 mag 2008 12:06:47 +0200

library ieee;
use ieee.std_logic_1164.all;

entity divisor is 
port (
    clk			: in	  std_logic); 
     
end divisor;     
        

architecture synth of divisor is
               
begin  

end synth;








